`timescale 1ns/1ps
import uvm_pkg::*;
`include "uvm_macros.svh"

`include "reg_model.sv"
`include "reg_block.sv"
`include "reg_seq_item.sv"
`include "reg_sequencer.sv"
`include "reg_interface.sv"
`include "reg_driver.sv"
`include "reg_sequence.sv" 
`include "reg_agent.sv"
`include "reg_adapter.sv"
`include "reg_env.sv"
`include "reg_test.sv"
`include "reg_design.sv"
`include "hdl_top.sv"
`include "hvl_top.sv"