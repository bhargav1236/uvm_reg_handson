module hvl_top;

import uvm_pkg::*;

initial begin
	run_test("reg_test");
end

endmodule